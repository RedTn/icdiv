magic
tech scmos
timestamp 1385276660
<< metal1 >>
rect -6 56 1 60
rect 9 42 11 46
rect 6 21 11 42
rect 102 17 105 31
rect -12 4 1 9
rect -12 -64 -6 4
rect -12 -68 0 -64
<< metal2 >>
rect -12 -12 -6 54
rect 95 42 105 46
rect 7 34 12 38
rect 93 34 100 38
rect -12 -17 -1 -12
rect 7 -28 11 17
rect 49 -8 53 10
rect 49 -11 61 -8
rect 7 -31 12 -28
rect 102 -35 105 12
rect 92 -39 105 -35
<< m2contact >>
rect -12 54 -6 60
rect 4 42 9 46
rect 100 31 105 38
rect 6 17 12 21
rect 102 12 106 17
rect -1 -18 3 -12
use 2to1muxfixed  2to1muxfixed_0
timestamp 1384797888
transform 1 0 31 0 1 35
box -31 -34 66 30
use 2to1muxfixed  2to1muxfixed_1
timestamp 1384797888
transform 1 0 31 0 1 -38
box -31 -34 66 30
<< end >>
