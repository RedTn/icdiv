magic
tech scmos
timestamp 1384799288
<< pwell >>
rect -12 -58 69 -28
<< nwell >>
rect -12 -28 69 4
<< polysilicon >>
rect 26 -3 30 -1
rect 46 -3 48 -1
rect 62 -3 64 -1
rect 26 -9 30 -7
rect -5 -11 -3 -9
rect 2 -11 4 -9
rect 46 -13 48 -7
rect 62 -8 64 -7
rect 54 -10 64 -8
rect 54 -15 56 -10
rect -5 -16 -3 -15
rect -7 -18 -3 -16
rect -7 -47 -5 -18
rect 2 -19 4 -15
rect 53 -17 56 -15
rect 15 -23 26 -19
rect 53 -20 55 -17
rect 2 -27 4 -23
rect 2 -31 6 -27
rect 49 -29 52 -22
rect 2 -47 4 -31
rect 49 -32 64 -29
rect 61 -33 64 -32
rect 42 -37 44 -36
rect 61 -39 64 -37
rect 30 -44 32 -42
rect 42 -43 44 -41
rect 18 -47 22 -44
rect 30 -46 40 -44
rect 38 -47 40 -46
rect -7 -53 -5 -51
rect 2 -53 4 -51
rect 18 -53 22 -51
rect 38 -53 40 -51
<< ndiffusion >>
rect 60 -37 61 -33
rect 64 -37 65 -33
rect 37 -41 42 -37
rect 44 -41 47 -37
rect -8 -51 -7 -47
rect -5 -51 -4 -47
rect 0 -51 2 -47
rect 4 -51 18 -47
rect 22 -51 25 -47
rect 37 -51 38 -47
rect 40 -51 47 -47
<< pdiffusion >>
rect 18 -7 26 -3
rect 30 -7 33 -3
rect 45 -7 46 -3
rect 48 -7 49 -3
rect 61 -7 62 -3
rect 64 -7 65 -3
rect -8 -15 -5 -11
rect -3 -15 2 -11
rect 4 -15 15 -11
rect 1 -23 2 -19
rect 4 -23 5 -19
<< metal1 >>
rect -20 0 -12 4
rect -4 0 77 4
rect -12 -11 -8 0
rect 14 -3 18 0
rect 41 -3 45 0
rect 57 -3 61 0
rect -1 -8 0 -5
rect -12 -19 -8 -15
rect -12 -23 -3 -19
rect 9 -23 11 -19
rect 10 -31 11 -27
rect 19 -35 23 -11
rect -12 -47 -8 -39
rect 19 -40 23 -39
rect 22 -44 23 -40
rect 26 -19 30 -13
rect 26 -40 30 -23
rect 33 -10 37 -7
rect 49 -10 53 -7
rect 33 -37 37 -14
rect 42 -19 46 -15
rect 49 -18 53 -14
rect 40 -32 44 -31
rect 65 -33 69 -7
rect 54 -37 55 -35
rect 26 -47 30 -44
rect 47 -47 51 -41
rect 29 -51 30 -47
rect -4 -54 0 -51
rect 33 -54 37 -51
rect 54 -54 58 -37
rect 65 -45 69 -37
rect -20 -58 55 -54
rect 65 -58 77 -54
<< metal2 >>
rect 29 0 33 8
rect 25 -4 33 0
rect 37 0 41 8
rect 37 -4 53 0
rect 4 -8 29 -4
rect 49 -10 53 -4
rect 37 -14 49 -10
rect 49 -19 53 -18
rect -20 -23 42 -19
rect 46 -23 77 -19
rect -20 -31 11 -27
rect 15 -31 40 -27
rect 44 -31 77 -27
rect -8 -39 19 -35
rect 29 -45 61 -41
rect 29 -62 33 -45
<< ntransistor >>
rect 61 -37 64 -33
rect 42 -41 44 -37
rect -7 -51 -5 -47
rect 2 -51 4 -47
rect 18 -51 22 -47
rect 38 -51 40 -47
<< ptransistor >>
rect 26 -7 30 -3
rect 46 -7 48 -3
rect 62 -7 64 -3
rect -5 -15 -3 -11
rect 2 -15 4 -11
rect 2 -23 4 -19
<< polycontact >>
rect -5 -9 -1 -5
rect 26 -13 30 -9
rect 42 -15 46 -11
rect 11 -23 15 -19
rect 26 -23 30 -19
rect 49 -22 53 -18
rect 6 -31 10 -27
rect 40 -36 44 -32
rect 18 -44 22 -40
rect 26 -44 30 -40
<< ndcontact >>
rect 55 -37 60 -33
rect 65 -37 69 -33
rect 33 -41 37 -37
rect 47 -41 51 -37
rect -12 -51 -8 -47
rect -4 -51 0 -47
rect 25 -51 29 -47
rect 33 -51 37 -47
rect 47 -51 51 -47
<< pdcontact >>
rect 14 -7 18 -3
rect 33 -7 37 -3
rect 41 -7 45 -3
rect 49 -7 53 -3
rect 57 -7 61 -3
rect 65 -7 69 -3
rect -12 -15 -8 -11
rect 15 -15 19 -11
rect -3 -23 1 -19
rect 5 -23 9 -19
<< m2contact >>
rect 0 -8 4 -4
rect 11 -31 15 -27
rect -12 -39 -8 -35
rect 19 -39 23 -35
rect 33 -14 37 -10
rect 42 -23 46 -19
rect 49 -14 53 -10
rect 40 -31 44 -27
rect 61 -45 65 -41
<< psubstratepcontact >>
rect 55 -58 65 -54
<< nsubstratencontact >>
rect -12 0 -4 4
<< labels >>
rlabel metal2 29 -4 33 8 1 D
rlabel metal2 29 -62 33 -41 5 Q
rlabel metal2 46 -23 77 -19 3 Rb
rlabel metal2 44 -31 77 -27 3 Clk
rlabel metal2 37 -4 41 8 1 Qb
<< end >>
