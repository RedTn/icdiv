magic
tech scmos
timestamp 1385773984
<< polysilicon >>
rect 63 -119 66 -113
rect 74 -118 77 -115
rect 84 -119 87 -115
<< metal1 >>
rect 151 87 282 88
rect -91 80 -8 84
rect -3 81 12 85
rect 91 81 282 87
rect -3 80 1 81
rect 130 80 263 81
rect 99 71 110 72
rect -91 68 4 71
rect -6 67 4 68
rect 103 67 281 71
rect -91 60 4 63
rect -6 59 4 60
rect 103 59 281 63
rect -6 58 8 59
rect 89 29 106 35
rect 113 29 232 35
rect 107 11 119 12
rect -3 6 10 10
rect 98 6 119 11
rect 98 -13 116 -12
rect -9 -14 3 -13
rect -94 -17 3 -14
rect 102 -17 281 -13
rect -9 -22 3 -21
rect -94 -25 3 -22
rect 102 -25 281 -21
rect -94 -26 8 -25
rect 99 -52 108 -47
rect 114 -52 231 -48
rect 93 -66 220 -65
rect 93 -72 207 -66
rect 206 -78 207 -72
rect 3 -94 119 -93
rect 11 -100 119 -94
rect 56 -113 62 -108
rect 74 -111 78 -108
rect 53 -114 67 -113
rect 83 -110 88 -104
rect 83 -111 93 -110
rect 87 -115 93 -111
rect 95 -122 119 -118
rect 104 -126 113 -125
rect 104 -127 108 -126
rect 101 -130 108 -127
rect 113 -130 232 -126
rect 17 -392 21 -357
rect 42 -371 45 -348
rect 68 -364 72 -338
rect 100 -345 126 -338
rect 111 -371 136 -370
rect 42 -375 136 -371
rect 17 -396 65 -392
rect 117 -419 152 -418
rect -94 -423 25 -419
rect 121 -423 281 -419
rect 133 -427 152 -426
rect -94 -431 15 -427
rect 117 -431 281 -427
rect 110 -461 126 -456
rect -54 -484 -19 -477
rect -84 -520 -9 -511
rect -5 -520 10 -511
rect -84 -521 10 -520
rect -27 -547 65 -543
rect 69 -547 70 -543
rect -27 -548 70 -547
rect -91 -596 35 -592
rect 41 -596 281 -592
rect -24 -606 44 -605
rect -91 -610 44 -606
rect 49 -606 238 -605
rect 49 -610 281 -606
rect -91 -611 281 -610
rect -13 -627 207 -623
rect -91 -639 179 -636
rect 185 -639 281 -636
rect -91 -650 191 -647
rect 196 -650 281 -647
rect -85 -718 -75 -712
rect 93 -829 128 -825
rect 132 -829 133 -825
rect 93 -830 133 -829
rect -91 -837 45 -833
rect 146 -837 281 -833
rect -91 -849 66 -845
rect 151 -849 281 -845
rect -91 -857 66 -853
rect 151 -857 281 -853
rect -91 -882 70 -881
rect -91 -886 66 -882
rect 151 -886 281 -882
rect -91 -894 66 -890
rect 146 -894 147 -890
rect 151 -894 281 -890
rect -91 -895 70 -894
rect 92 -910 97 -907
rect 96 -915 97 -910
rect -77 -945 -76 -939
rect -71 -945 54 -939
rect -90 -966 51 -962
rect 148 -966 281 -962
rect -90 -974 51 -970
rect 148 -974 281 -970
rect -88 -1002 -55 -998
rect -48 -1003 53 -997
rect 147 -1003 230 -996
rect 237 -1003 280 -996
rect 99 -1016 100 -1012
rect 104 -1016 207 -1012
<< metal2 >>
rect 55 85 59 90
rect -8 10 -3 80
rect 54 12 58 34
rect 63 21 67 29
rect 62 12 67 21
rect -8 6 -7 10
rect 107 -47 113 29
rect 107 -52 108 -47
rect 54 -57 78 -53
rect -77 -484 -61 -477
rect -89 -712 -85 -522
rect -77 -541 -73 -484
rect -78 -581 -73 -541
rect -34 -543 -27 -83
rect 2 -94 11 -93
rect 2 -116 11 -100
rect 50 -108 55 -81
rect 74 -104 78 -57
rect 88 -104 93 -72
rect 2 -263 10 -116
rect 108 -126 114 -52
rect 119 -93 124 6
rect 232 -46 236 29
rect 119 -118 124 -100
rect 123 -122 124 -118
rect 113 -130 114 -126
rect 3 -412 10 -263
rect 208 -286 218 -78
rect 207 -296 218 -286
rect 232 -126 236 -52
rect 72 -368 77 -364
rect 65 -403 69 -396
rect 73 -404 77 -368
rect 126 -455 132 -345
rect 130 -460 132 -455
rect -13 -484 18 -477
rect -78 -666 -74 -581
rect -17 -650 -13 -627
rect -9 -650 -5 -520
rect 65 -543 69 -536
rect 136 -546 140 -375
rect 65 -556 69 -547
rect 73 -550 140 -546
rect 73 -555 77 -550
rect 35 -654 39 -597
rect 44 -654 48 -610
rect 136 -652 140 -550
rect 207 -623 217 -296
rect 216 -627 217 -623
rect 207 -629 217 -627
rect 179 -657 185 -640
rect 207 -655 216 -629
rect -76 -939 -71 -733
rect -54 -997 -49 -789
rect 129 -807 133 -805
rect 127 -809 133 -807
rect 46 -814 133 -809
rect 46 -832 51 -814
rect 129 -825 133 -814
rect 132 -829 133 -825
rect 96 -915 104 -910
rect 100 -937 104 -915
rect 100 -1011 104 -1002
rect 207 -1012 215 -655
rect 232 -996 236 -130
<< polycontact >>
rect 62 -113 67 -108
rect 73 -115 78 -111
rect 83 -115 87 -111
<< m2contact >>
rect -8 80 -3 85
rect 4 67 8 71
rect 99 67 103 71
rect 4 59 8 63
rect 97 59 103 63
rect 106 29 113 35
rect 232 29 238 35
rect -7 6 -3 10
rect 119 6 125 12
rect 3 -17 8 -13
rect 98 -17 102 -13
rect 3 -25 8 -21
rect 98 -25 102 -21
rect 108 -52 114 -47
rect 231 -52 238 -46
rect 88 -72 93 -65
rect 207 -78 220 -66
rect 2 -100 11 -94
rect 119 -100 125 -93
rect 74 -108 78 -104
rect 50 -113 56 -108
rect 88 -110 93 -104
rect 119 -122 123 -118
rect 108 -130 113 -126
rect 232 -130 236 -126
rect 126 -345 133 -338
rect 68 -368 72 -364
rect 136 -375 140 -370
rect 65 -396 69 -392
rect 117 -423 121 -419
rect 15 -431 19 -427
rect 126 -461 130 -455
rect -61 -484 -54 -477
rect -19 -484 -13 -477
rect -89 -522 -84 -511
rect -9 -520 -5 -511
rect -34 -549 -27 -543
rect 65 -547 69 -543
rect 35 -597 41 -591
rect 44 -610 49 -605
rect -17 -627 -13 -623
rect 207 -627 216 -623
rect 179 -640 185 -635
rect 191 -654 196 -645
rect -89 -718 -85 -712
rect -54 -789 -48 -785
rect 128 -829 132 -825
rect 45 -837 52 -832
rect 66 -849 70 -845
rect 147 -849 151 -845
rect 66 -857 70 -853
rect 147 -857 151 -853
rect 66 -886 70 -882
rect 147 -886 151 -882
rect 66 -894 70 -890
rect 147 -894 151 -890
rect 92 -915 96 -910
rect -76 -945 -71 -939
rect 51 -966 55 -962
rect 144 -966 148 -962
rect 51 -974 55 -970
rect 144 -974 148 -970
rect -55 -1004 -48 -997
rect 230 -1003 237 -996
rect 100 -1016 104 -1011
rect 207 -1017 216 -1012
use 2to1mux  2to1mux_0
timestamp 1384565173
transform 1 0 37 0 1 60
box -31 -34 66 30
use dflipfloplabels  dflipfloplabels_0
timestamp 1384799288
transform 1 0 25 0 1 6
box -20 -62 77 8
use addsub1  addsub1_0
timestamp 1385343589
transform 1 0 77 0 1 -139
box -74 -223 37 25
use real21mux  real21mux_0
timestamp 1385276660
transform 1 0 16 0 1 -465
box -12 -72 106 65
use real31mux  real31mux_0
timestamp 1385664840
transform 1 0 -84 0 1 -793
box 6 -14 280 146
use shiftv2  shiftv2_0
timestamp 1385333955
transform 1 0 101 0 1 -902
box -35 -8 50 73
use dflipfloplabels  dflipfloplabels_1
timestamp 1384799288
transform 1 0 71 0 1 -943
box -20 -62 77 8
<< labels >>
rlabel metal2 65 -555 69 -552 1 c
rlabel metal1 91 81 132 87 1 Vdd
rlabel metal2 74 -85 77 -83 1 b
rlabel metal1 156 -430 166 -427 1 add
rlabel metal1 141 -422 155 -422 1 addb
rlabel metal2 73 -555 77 -552 1 a
rlabel metal2 88 -83 92 -81 1 aa
rlabel metal2 51 -87 54 -83 1 cc
rlabel space -22 -1004 10 -997 1 GND
rlabel metal2 232 -920 236 -917 1 GND
rlabel metal1 171 59 179 63 1 l
rlabel metal1 202 -17 210 -13 1 tb
rlabel metal2 55 85 59 90 1 in
rlabel metal1 189 -24 192 -22 1 clk
rlabel metal1 186 69 190 70 1 lb
rlabel metal2 63 16 66 20 1 bb
rlabel metal2 54 16 57 20 1 out
<< end >>
