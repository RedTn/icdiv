magic
tech scmos
timestamp 1384797888
<< pwell >>
rect -9 -30 47 -5
<< nwell >>
rect -9 -5 47 25
<< polysilicon >>
rect 12 11 14 13
rect 23 11 25 13
rect 31 11 33 13
rect 39 11 41 13
rect -4 4 -2 6
rect 12 3 14 7
rect -4 -10 -2 0
rect 12 -3 14 -1
rect 7 -5 14 -3
rect 12 -7 14 -5
rect 12 -9 17 -7
rect 15 -10 17 -9
rect 23 -10 25 7
rect -4 -16 -2 -14
rect 15 -16 17 -14
rect 23 -16 25 -14
rect 31 -18 33 7
rect 39 4 41 7
rect 39 2 42 4
rect 40 -9 42 2
rect 39 -12 42 -9
rect 39 -18 41 -12
rect 31 -24 33 -22
rect 39 -24 41 -22
<< ndiffusion >>
rect -5 -14 -4 -10
rect -2 -14 -1 -10
rect 14 -14 15 -10
rect 17 -14 18 -10
rect 22 -14 23 -10
rect 25 -14 26 -10
rect 30 -22 31 -18
rect 33 -22 34 -18
rect 38 -22 39 -18
rect 41 -22 42 -18
<< pdiffusion >>
rect 11 7 12 11
rect 14 7 23 11
rect 25 7 26 11
rect 30 7 31 11
rect 33 7 39 11
rect 41 7 43 11
rect -5 0 -4 4
rect -2 0 -1 4
<< metal1 >>
rect -31 21 -9 25
rect 47 21 66 25
rect -16 -3 -12 14
rect -9 11 -5 21
rect -9 7 7 11
rect 18 8 22 12
rect 43 11 47 21
rect -9 4 -5 7
rect 3 -2 7 4
rect 19 3 22 8
rect -16 -7 -8 -3
rect 26 -4 30 7
rect 52 0 56 14
rect 34 -2 38 -1
rect 19 -5 30 -4
rect 3 -14 7 -6
rect 22 -7 30 -5
rect 46 -4 56 0
rect 18 -10 22 -9
rect 52 -9 56 -4
rect 30 -14 46 -10
rect -9 -26 -5 -14
rect 11 -18 14 -14
rect 26 -18 30 -14
rect 42 -18 46 -14
rect 11 -22 26 -18
rect 34 -26 38 -22
rect -31 -30 -9 -26
rect 22 -30 66 -26
<< metal2 >>
rect 18 24 22 30
rect 10 20 22 24
rect 26 22 30 30
rect 10 19 14 20
rect -16 18 14 19
rect 26 18 56 22
rect -12 15 14 18
rect 18 11 22 12
rect -31 10 -20 11
rect -8 10 48 11
rect 60 10 66 11
rect -31 7 66 10
rect -31 -1 34 3
rect 38 -1 66 3
rect 18 -34 22 -9
rect 36 -13 52 -9
rect 36 -26 40 -13
rect 44 -14 47 -13
rect 26 -30 40 -26
rect 26 -34 30 -30
<< ntransistor >>
rect -4 -14 -2 -10
rect 15 -14 17 -10
rect 23 -14 25 -10
rect 31 -22 33 -18
rect 39 -22 41 -18
<< ptransistor >>
rect 12 7 14 11
rect 23 7 25 11
rect 31 7 33 11
rect 39 7 41 11
rect -4 0 -2 4
<< polycontact >>
rect -8 -7 -4 -3
rect 12 -1 16 3
rect 19 -1 23 3
rect 3 -6 7 -2
rect 33 -6 37 -2
rect 42 -4 46 0
<< ndcontact >>
rect -9 -14 -5 -10
rect -1 -14 3 -10
rect 10 -14 14 -10
rect 18 -14 22 -10
rect 26 -14 30 -10
rect 26 -22 30 -18
rect 34 -22 38 -18
rect 42 -22 46 -18
<< pdcontact >>
rect 7 7 11 11
rect 26 7 30 11
rect 43 7 47 11
rect -9 0 -5 4
rect -1 0 3 4
<< m2contact >>
rect -16 14 -12 18
rect 18 12 22 16
rect 52 14 56 18
rect 34 -1 38 3
rect 18 -9 22 -5
rect 52 -13 56 -9
<< psubstratepcontact >>
rect -9 -30 22 -26
<< nsubstratencontact >>
rect -9 21 47 25
<< labels >>
rlabel nwell -9 -5 47 25 8 Vdd
rlabel pwell -9 -30 47 -5 6 Gnd
rlabel metal2 26 -34 30 -26 5 Qb
rlabel metal2 18 -34 22 -9 5 D
rlabel metal2 18 20 22 30 1 divisor
rlabel space -8 7 58 11 3 loadb
rlabel metal2 38 -1 58 3 3 load
<< end >>
