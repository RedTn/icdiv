magic
tech scmos
timestamp 1385774014
<< metal1 >>
rect 6188 1277 7380 1282
rect 6318 1238 6319 1250
rect 6334 1238 7314 1250
rect 6318 1237 7314 1238
rect 6352 1211 6856 1216
rect 6851 1100 6856 1211
rect 6855 1096 6856 1100
rect 667 1075 676 1083
rect 3111 1078 5925 1085
rect 6770 1074 6787 1078
rect 3122 1064 6584 1068
rect 3120 1056 6594 1060
rect 392 1028 413 1032
rect 3112 980 6347 984
rect 3104 972 6444 976
rect 463 910 725 915
rect 735 910 736 915
rect 817 910 1059 915
rect 1151 911 1392 915
rect 1483 910 1742 914
rect 1833 911 2102 915
rect 2192 911 2327 917
rect 2382 911 2449 917
rect 2321 905 2388 911
rect 2540 909 2805 915
rect 2881 917 2886 948
rect 6851 940 6856 1096
rect 6981 1131 7233 1135
rect 6710 897 6715 935
rect 6538 829 6612 833
rect 6509 817 6610 818
rect 6513 813 6609 817
rect 6487 798 6591 801
rect 6384 781 6599 785
rect 6384 780 6603 781
rect 6238 749 6611 753
rect 6414 733 6599 737
rect 6288 725 6610 729
rect 6981 705 6985 1131
rect 7301 1119 7314 1237
rect 6800 701 6985 705
rect 2971 651 3011 655
rect 3007 627 3011 651
rect 3007 623 6177 627
rect 6188 623 6426 627
rect 6432 623 6609 627
rect 5932 607 6320 611
rect 6332 607 6460 611
rect 6464 607 6612 611
rect 3120 574 6371 578
rect 3118 566 6401 570
rect 3016 459 6564 470
rect 3017 430 3028 459
rect 548 421 3028 430
rect 3118 425 3175 430
rect 3118 401 3123 425
rect 6094 424 6524 428
rect 3134 412 3180 416
rect 3134 392 3140 412
rect 6049 410 6497 414
rect 3149 398 3159 399
rect 3117 385 3140 392
rect 3148 393 3176 398
rect 3148 392 3159 393
rect 6050 392 6590 396
rect 3148 362 3154 392
rect 3122 357 3154 362
rect 3161 379 3176 383
rect 3161 350 3166 379
rect 6096 377 6552 381
rect 3121 347 3166 350
rect 937 330 1023 339
rect 3015 337 3159 338
rect 3173 337 3188 345
rect 6113 341 6481 345
rect 3015 331 3188 337
rect 6096 327 6100 341
rect 6096 323 6459 327
rect 932 208 1020 216
rect 6107 174 6111 285
rect 3119 169 3178 173
rect 6097 170 6111 174
rect 3119 164 3123 169
rect 6100 167 6108 170
rect 3131 157 3176 161
rect 3131 152 3138 157
rect 6098 155 6233 159
rect 3119 148 3138 152
rect 3174 144 3178 153
rect 6081 147 6282 151
rect 3122 140 3178 144
rect 3121 120 3177 124
rect 3121 111 3125 120
rect 6097 118 6282 122
rect 3168 107 3177 115
rect 6094 110 6231 114
rect 3118 103 3177 107
rect 910 54 1022 58
rect 3118 40 3176 44
rect 3118 31 3126 40
rect 6099 38 6349 42
rect 3173 27 3178 35
rect 6097 30 6441 34
rect 6449 30 6863 34
rect 3121 23 3178 27
rect 1034 -9 1057 4
rect 3112 -5 3182 9
rect 6097 3 6426 7
rect 7375 -97 7380 1277
rect 7282 -101 7380 -97
<< metal2 >>
rect 6177 1282 6188 1306
rect 387 1090 466 1094
rect 387 1032 391 1090
rect 462 1086 466 1090
rect 817 1085 821 1161
rect 1149 1086 1153 1161
rect 1482 1086 1486 1161
rect 1832 1086 1836 1161
rect 2192 1086 2196 1161
rect 2540 1085 2544 1161
rect 2897 1085 2901 1161
rect 2559 926 2563 929
rect 2886 913 2898 916
rect 3269 534 3274 1161
rect 3635 535 3640 1161
rect 4001 535 4006 1161
rect 3269 519 3275 534
rect 3635 520 3641 535
rect 4001 520 4007 535
rect 3269 510 3274 519
rect 4001 518 4006 520
rect 4367 519 4373 1161
rect 4731 536 4736 1161
rect 4731 520 4737 536
rect 4731 515 4736 520
rect 5098 517 5104 1161
rect 5461 534 5466 1161
rect 5825 534 5830 1161
rect 5928 611 5932 1078
rect 6177 627 6188 1276
rect 6320 1251 6333 1303
rect 6233 749 6234 753
rect 5461 518 5467 534
rect 5825 518 5831 534
rect 5461 508 5466 518
rect 5825 494 5830 518
rect 2622 453 2625 458
rect 6106 289 6110 341
rect 6106 285 6107 289
rect 3404 187 3410 192
rect 6233 160 6238 749
rect 6233 114 6238 155
rect 6283 152 6287 725
rect 6320 611 6333 1238
rect 6348 999 6352 1211
rect 6805 1102 6809 1354
rect 6778 1098 6818 1102
rect 6757 1074 6770 1078
rect 6835 1078 6839 1352
rect 7234 1135 7238 1341
rect 7234 1126 7238 1130
rect 6855 1096 7185 1100
rect 6794 1074 7172 1078
rect 6348 986 6353 999
rect 6332 606 6333 611
rect 6283 123 6287 146
rect 6349 42 6353 980
rect 6442 972 6444 976
rect 6448 972 6449 976
rect 6372 580 6382 779
rect 6403 574 6413 732
rect 6426 12 6432 623
rect 6442 35 6449 972
rect 6529 829 6532 833
rect 6500 813 6509 817
rect 6513 813 6514 817
rect 6481 797 6482 801
rect 6460 327 6464 607
rect 6481 347 6487 797
rect 6500 415 6504 813
rect 6529 795 6533 829
rect 6585 809 6588 1064
rect 6595 848 6600 1056
rect 6715 935 6851 940
rect 6596 825 6600 848
rect 6611 829 6612 833
rect 6617 829 6619 833
rect 6596 821 6623 825
rect 6613 813 6620 817
rect 6585 805 6621 809
rect 6595 798 6619 801
rect 6526 791 6533 795
rect 6526 431 6530 791
rect 6553 789 6619 793
rect 6553 382 6557 789
rect 6604 781 6622 785
rect 6615 749 6619 753
rect 6603 733 6623 737
rect 6614 725 6623 729
rect 6725 701 6794 705
rect 6567 676 6619 680
rect 6567 470 6575 676
rect 6613 623 6619 627
rect 6592 615 6619 619
rect 6592 397 6596 615
rect 6616 607 6619 611
rect 6460 322 6464 323
rect 6863 34 6867 1074
rect 507 -151 511 -16
rect 862 -151 866 -15
rect 1194 -151 1198 -16
rect 1527 -151 1531 -16
rect 1877 -151 1881 -16
rect 2237 -151 2241 -15
rect 2585 -151 2589 -16
rect 2942 -151 2946 -17
rect 3395 -151 3399 -5
rect 3761 -151 3765 -5
rect 4127 -151 4131 -4
rect 4493 -151 4497 -2
rect 4857 -151 4861 -6
rect 5224 -151 5228 -6
rect 5587 -151 5591 -6
rect 5951 -151 5955 -6
rect 7234 -119 7238 -93
<< m2contact >>
rect 6176 1276 6188 1282
rect 6319 1238 6334 1251
rect 6348 1211 6352 1216
rect 6851 1096 6855 1100
rect 5925 1078 5936 1093
rect 6787 1071 6794 1080
rect 6584 1064 6589 1069
rect 6594 1056 6601 1061
rect 386 1028 392 1032
rect 6347 980 6353 986
rect 6444 972 6448 976
rect 455 909 463 920
rect 725 908 735 915
rect 808 907 817 918
rect 1059 908 1069 916
rect 1142 908 1151 918
rect 1392 910 1401 916
rect 1476 909 1483 916
rect 1742 908 1751 915
rect 1826 910 1833 916
rect 2102 910 2111 916
rect 2185 909 2192 918
rect 2449 909 2460 918
rect 2533 909 2540 917
rect 2805 907 2816 918
rect 2880 912 2886 917
rect 6710 935 6715 940
rect 6851 935 6856 940
rect 6710 892 6715 897
rect 6532 829 6538 833
rect 6612 829 6617 833
rect 6509 813 6513 817
rect 6609 813 6613 817
rect 6482 797 6487 801
rect 6591 797 6595 801
rect 6372 779 6384 786
rect 6599 781 6604 785
rect 6234 749 6238 753
rect 6611 749 6615 753
rect 6403 732 6414 741
rect 6599 733 6603 737
rect 6283 725 6288 730
rect 6610 725 6614 729
rect 7233 1130 7238 1135
rect 6794 701 6800 705
rect 6177 623 6188 627
rect 6426 623 6432 627
rect 6609 623 6613 627
rect 5928 607 5932 611
rect 6320 606 6332 611
rect 6460 607 6464 611
rect 6612 607 6616 611
rect 6371 574 6382 580
rect 6401 566 6415 574
rect 6564 459 6575 470
rect 542 420 548 432
rect 6524 421 6533 431
rect 6497 408 6506 415
rect 6590 392 6597 397
rect 6552 377 6557 382
rect 6106 341 6113 346
rect 6481 341 6487 347
rect 6459 323 6465 327
rect 6107 285 6111 289
rect 6233 155 6238 160
rect 6282 146 6287 152
rect 6282 118 6288 123
rect 6231 109 6239 114
rect 6349 38 6353 42
rect 6441 29 6449 35
rect 6863 30 6867 34
rect 6426 3 6432 12
use highdata  highdata_1
timestamp 1385774014
transform 1 0 407 0 1 998
box -94 -1017 282 90
use highdata  highdata_2
timestamp 1385774014
transform 1 0 762 0 1 997
box -94 -1017 282 90
use highdata  highdata_3
timestamp 1385774014
transform 1 0 1094 0 1 997
box -94 -1017 282 90
use highdata  highdata_4
timestamp 1385774014
transform 1 0 1427 0 1 997
box -94 -1017 282 90
use highdata  highdata_5
timestamp 1385774014
transform 1 0 1777 0 1 997
box -94 -1017 282 90
use highdata  highdata_6
timestamp 1385774014
transform 1 0 2137 0 1 997
box -94 -1017 282 90
use highdata  highdata_7
timestamp 1385774014
transform 1 0 2485 0 1 997
box -94 -1017 282 90
use highdata  highdata_8
timestamp 1385774014
transform 1 0 2842 0 1 997
box -94 -1017 282 90
use controller_v2  controller_v2_0
timestamp 1384924723
transform 0 1 6661 -1 0 1079
box -105 -42 472 132
use lowdata  lowdata_0
timestamp 1385774014
transform 1 0 3203 0 1 206
box -29 -216 341 319
use lowdata  lowdata_1
timestamp 1385774014
transform 1 0 3569 0 1 206
box -29 -216 341 319
use lowdata  lowdata_2
timestamp 1385774014
transform 1 0 3935 0 1 206
box -29 -216 341 319
use lowdata  lowdata_3
timestamp 1385774014
transform 1 0 4301 0 1 206
box -29 -216 341 319
use lowdata  lowdata_4
timestamp 1385774014
transform 1 0 4665 0 1 205
box -29 -216 341 319
use lowdata  lowdata_5
timestamp 1385774014
transform 1 0 5032 0 1 205
box -29 -216 341 319
use lowdata  lowdata_6
timestamp 1385774014
transform 1 0 5395 0 1 204
box -29 -216 341 319
use lowdata  lowdata_7
timestamp 1385774014
transform 1 0 5759 0 1 204
box -29 -216 341 319
use value  value_0
timestamp 1385683202
transform 1 0 7185 0 1 1057
box -35 -1162 135 70
<< labels >>
rlabel metal1 6581 623 6587 626 1 GND
rlabel metal1 6580 607 6584 611 1 Vdd
rlabel metal2 6788 702 6798 705 1 start
rlabel metal1 6588 749 6596 753 1 shift
rlabel metal2 2622 453 2625 458 1 testt
rlabel metal2 6598 845 6600 850 1 test3
rlabel metal2 6824 1074 6837 1078 1 clk
rlabel metal1 3000 652 3011 654 1 GND
rlabel space 6084 341 6090 345 1 Vdd
rlabel metal1 6556 799 6559 801 1 inbit
rlabel metal1 6397 378 6401 381 1 sel0
rlabel metal1 6405 411 6407 413 1 sel1
rlabel metal1 3447 980 3455 983 1 rstb
rlabel metal2 2897 1147 2901 1160 1 divisorin_0
rlabel metal2 2541 1149 2544 1160 1 divisorin_1
rlabel metal2 2192 1149 2196 1161 1 divisorin_2
rlabel metal2 1833 1147 1836 1160 1 divisorin_3
rlabel metal2 1483 1147 1486 1160 1 divisorin_4
rlabel metal2 1149 1146 1153 1157 1 divisorin_5
rlabel metal2 817 1147 821 1159 1 divisorin_6
rlabel metal2 5826 1147 5829 1157 1 dividendin_0
rlabel metal2 5462 1146 5465 1159 1 dividendin_1
rlabel metal2 5099 1147 5102 1160 1 dividendin_2
rlabel metal2 4733 1147 4736 1160 1 dividendin_3
rlabel metal2 4367 1147 4370 1160 1 dividendin_4
rlabel metal2 4001 1146 4004 1159 1 dividendin_5
rlabel metal2 3636 1148 3639 1161 1 dividendin_6
rlabel metal2 3270 1146 3273 1159 1 dividendin_7
rlabel metal2 5952 -146 5955 -132 1 quotient_0
rlabel metal2 5588 -143 5591 -129 1 quotient_1
rlabel metal2 5225 -141 5228 -127 1 quotient_2
rlabel metal2 4857 -146 4860 -132 1 quotient_3
rlabel metal2 4494 -142 4497 -128 1 quotient_4
rlabel metal2 4128 -141 4131 -127 1 quotient_5
rlabel metal2 3762 -143 3765 -129 1 quotient_6
rlabel metal2 3396 -139 3399 -125 1 quotient_7
rlabel metal2 2585 -145 2588 -134 1 remainder_0
rlabel metal2 2238 -141 2241 -132 1 remainder_1
rlabel metal2 1877 -143 1880 -134 1 remainder_2
rlabel metal2 1528 -142 1531 -133 1 remainder_3
rlabel metal2 1195 -140 1198 -131 1 remainder_4
rlabel metal2 863 -144 866 -135 1 remainder_5
rlabel metal2 508 -148 511 -139 1 remainder_6
rlabel metal2 6807 1119 6808 1124 1 reset
rlabel metal2 7236 -117 7237 -110 1 value
<< end >>
