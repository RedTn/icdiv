magic
tech scmos
timestamp 1385698489
<< metal1 >>
rect 667 1075 676 1083
rect 3111 1078 3148 1085
rect 3122 1064 3148 1068
rect 3120 1056 3148 1060
rect 392 1028 413 1032
rect 3112 980 3148 984
rect 3104 972 3148 976
rect 463 910 725 915
rect 735 910 736 915
rect 817 910 1059 915
rect 1151 911 1392 915
rect 1483 910 1742 914
rect 1833 911 2102 915
rect 2192 911 2327 917
rect 2382 911 2449 917
rect 2321 905 2388 911
rect 2540 909 2805 915
rect 2881 917 2886 948
rect 2971 651 3011 655
rect 3007 627 3011 651
rect 3007 623 3148 627
rect 3120 574 3148 578
rect 3118 566 3148 570
rect 3016 459 6138 470
rect 3017 430 3028 459
rect 548 421 3028 430
rect 3118 425 3175 430
rect 3118 401 3123 425
rect 6094 424 6148 428
rect 3134 412 3180 416
rect 3134 392 3140 412
rect 6049 410 6145 414
rect 3149 398 3159 399
rect 3117 385 3140 392
rect 3148 393 3176 398
rect 3148 392 3159 393
rect 6050 392 6148 396
rect 3148 362 3154 392
rect 3122 357 3154 362
rect 3161 379 3176 383
rect 3161 350 3166 379
rect 6096 377 6148 381
rect 3121 347 3166 350
rect 937 330 1023 339
rect 3015 337 3159 338
rect 3173 337 3188 345
rect 3015 331 3188 337
rect 932 208 1020 216
rect 6107 174 6111 224
rect 3119 169 3178 173
rect 6097 170 6111 174
rect 3119 164 3123 169
rect 6100 167 6108 170
rect 3131 157 3176 161
rect 3131 152 3138 157
rect 6098 155 6138 159
rect 3119 148 3138 152
rect 3174 144 3178 153
rect 6081 147 6138 151
rect 3122 140 3178 144
rect 3121 120 3177 124
rect 3121 111 3125 120
rect 6097 118 6138 122
rect 3168 107 3177 115
rect 6094 110 6138 114
rect 3118 103 3177 107
rect 910 54 1022 58
rect 3118 40 3176 44
rect 3118 31 3126 40
rect 6099 38 6138 42
rect 3173 27 3178 35
rect 6097 30 6138 34
rect 3121 23 3178 27
rect 1034 -9 1057 4
rect 3112 -5 3182 9
rect 6097 3 6138 7
<< metal2 >>
rect 387 1090 466 1094
rect 387 1032 391 1090
rect 462 1086 466 1090
rect 817 1085 821 1161
rect 1149 1086 1153 1161
rect 1482 1086 1486 1161
rect 1832 1086 1836 1161
rect 2192 1086 2196 1161
rect 2540 1085 2544 1161
rect 2897 1085 2901 1161
rect 2559 926 2563 929
rect 2886 913 2898 916
rect 3269 534 3274 1161
rect 3635 535 3640 1161
rect 4001 535 4006 1161
rect 3269 519 3275 534
rect 3635 520 3641 535
rect 4001 520 4007 535
rect 3269 510 3274 519
rect 4001 518 4006 520
rect 4367 519 4373 1161
rect 4731 536 4736 1161
rect 4731 520 4737 536
rect 4731 515 4736 520
rect 5098 517 5104 1161
rect 5461 534 5466 1161
rect 5825 534 5830 1161
rect 5461 518 5467 534
rect 5825 518 5831 534
rect 5461 508 5466 518
rect 5825 494 5830 518
rect 2622 453 2625 458
rect 3404 187 3410 192
rect 507 -151 511 -16
rect 862 -151 866 -15
rect 1194 -151 1198 -16
rect 1527 -151 1531 -16
rect 1877 -151 1881 -16
rect 2237 -151 2241 -15
rect 2585 -151 2589 -16
rect 2942 -151 2946 -17
rect 3395 -151 3399 -5
rect 3761 -151 3765 -5
rect 4127 -151 4131 -4
rect 4493 -151 4497 -2
rect 4857 -151 4861 -6
rect 5224 -151 5228 -6
rect 5587 -151 5591 -6
rect 5951 -151 5955 -6
<< m2contact >>
rect 386 1028 392 1032
rect 455 909 463 920
rect 725 908 735 915
rect 808 907 817 918
rect 1059 908 1069 916
rect 1142 908 1151 918
rect 1392 910 1401 916
rect 1476 909 1483 916
rect 1742 908 1751 915
rect 1826 910 1833 916
rect 2102 910 2111 916
rect 2185 909 2192 918
rect 2449 909 2460 918
rect 2533 909 2540 917
rect 2805 907 2816 918
rect 2880 912 2886 917
rect 542 420 548 432
use highdata  highdata_1
timestamp 1385698489
transform 1 0 407 0 1 998
box -94 -1017 282 90
use highdata  highdata_2
timestamp 1385698489
transform 1 0 762 0 1 997
box -94 -1017 282 90
use highdata  highdata_3
timestamp 1385698489
transform 1 0 1094 0 1 997
box -94 -1017 282 90
use highdata  highdata_4
timestamp 1385698489
transform 1 0 1427 0 1 997
box -94 -1017 282 90
use highdata  highdata_5
timestamp 1385698489
transform 1 0 1777 0 1 997
box -94 -1017 282 90
use highdata  highdata_6
timestamp 1385698489
transform 1 0 2137 0 1 997
box -94 -1017 282 90
use highdata  highdata_7
timestamp 1385698489
transform 1 0 2485 0 1 997
box -94 -1017 282 90
use highdata  highdata_8
timestamp 1385698489
transform 1 0 2842 0 1 997
box -94 -1017 282 90
use lowdata  lowdata_0
timestamp 1385698489
transform 1 0 3203 0 1 206
box -29 -216 341 319
use lowdata  lowdata_1
timestamp 1385698489
transform 1 0 3569 0 1 206
box -29 -216 341 319
use lowdata  lowdata_2
timestamp 1385698489
transform 1 0 3935 0 1 206
box -29 -216 341 319
use lowdata  lowdata_3
timestamp 1385698489
transform 1 0 4301 0 1 206
box -29 -216 341 319
use lowdata  lowdata_4
timestamp 1385698489
transform 1 0 4665 0 1 205
box -29 -216 341 319
use lowdata  lowdata_5
timestamp 1385698489
transform 1 0 5032 0 1 205
box -29 -216 341 319
use lowdata  lowdata_6
timestamp 1385698489
transform 1 0 5395 0 1 204
box -29 -216 341 319
use lowdata  lowdata_7
timestamp 1385698489
transform 1 0 5759 0 1 204
box -29 -216 341 319
<< labels >>
rlabel metal2 2622 453 2625 458 1 testt
rlabel metal1 3000 652 3011 654 1 GND
rlabel space 6084 341 6090 345 1 Vdd
rlabel metal2 2897 1147 2901 1160 1 divisorin_0
rlabel metal2 2541 1149 2544 1160 1 divisorin_1
rlabel metal2 2192 1149 2196 1161 1 divisorin_2
rlabel metal2 1833 1147 1836 1160 1 divisorin_3
rlabel metal2 1483 1147 1486 1160 1 divisorin_4
rlabel metal2 1149 1146 1153 1157 1 divisorin_5
rlabel metal2 817 1147 821 1159 1 divisorin_6
rlabel metal2 5826 1147 5829 1157 1 dividendin_0
rlabel metal2 5462 1146 5465 1159 1 dividendin_1
rlabel metal2 5099 1147 5102 1160 1 dividendin_2
rlabel metal2 4733 1147 4736 1160 1 dividendin_3
rlabel metal2 4367 1147 4370 1160 1 dividendin_4
rlabel metal2 4001 1146 4004 1159 1 dividendin_5
rlabel metal2 3636 1148 3639 1161 1 dividendin_6
rlabel metal2 3270 1146 3273 1159 1 dividendin_7
rlabel metal2 5952 -146 5955 -132 1 quotient_0
rlabel metal2 5588 -143 5591 -129 1 quotient_1
rlabel metal2 5225 -141 5228 -127 1 quotient_2
rlabel metal2 4857 -146 4860 -132 1 quotient_3
rlabel metal2 4494 -142 4497 -128 1 quotient_4
rlabel metal2 4128 -141 4131 -127 1 quotient_5
rlabel metal2 3762 -143 3765 -129 1 quotient_6
rlabel metal2 3396 -139 3399 -125 1 quotient_7
rlabel metal2 2585 -145 2588 -134 1 remainder_0
rlabel metal2 2238 -141 2241 -132 1 remainder_1
rlabel metal2 1877 -143 1880 -134 1 remainder_2
rlabel metal2 1528 -142 1531 -133 1 remainder_3
rlabel metal2 1195 -140 1198 -131 1 remainder_4
rlabel metal2 863 -144 866 -135 1 remainder_5
rlabel metal2 508 -148 511 -139 1 remainder_6
rlabel metal1 6110 148 6114 151 1 shiftb
rlabel metal1 6108 186 6110 190 1 inbit
rlabel metal1 6114 156 6121 158 1 shift
rlabel metal1 6119 120 6122 122 1 shiftb
rlabel metal1 6113 111 6120 113 1 shift
rlabel metal1 3136 624 3142 627 1 GND
rlabel metal1 3136 577 3139 577 1 addb
rlabel metal1 3136 567 3139 569 1 add
rlabel metal1 6126 39 6134 42 1 resetb
rlabel metal1 6125 31 6129 33 1 clk
rlabel metal1 3137 1065 3141 1067 1 loadb
rlabel metal1 3137 1057 3140 1058 1 load
rlabel metal1 3136 981 3139 983 1 resetb
rlabel metal1 3141 974 3144 975 1 clk
rlabel metal1 3129 1083 3139 1084 1 Vdd
rlabel metal1 6142 379 6146 380 7 sel_1
rlabel metal1 6139 393 6143 394 1 selb_1
rlabel metal1 6140 412 6144 413 1 sel_0
rlabel metal1 6139 425 6146 427 1 selb_0
<< end >>
