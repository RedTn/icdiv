magic
tech scmos
timestamp 1384720590
<< pwell >>
rect -10 -18 18 -3
<< nwell >>
rect -10 -3 18 12
<< polysilicon >>
rect -1 6 1 9
rect -1 0 1 2
rect 7 -8 9 -6
rect 7 -15 9 -12
<< ndiffusion >>
rect 6 -12 7 -8
rect 9 -12 10 -8
<< pdiffusion >>
rect -2 2 -1 6
rect 1 2 2 6
<< metal1 >>
rect -2 13 2 14
rect 6 2 14 6
rect -6 -1 -2 2
rect -10 -5 -2 -1
rect -6 -8 -2 -5
rect 10 -1 14 2
rect 10 -5 18 -1
rect 10 -8 14 -5
rect -6 -12 2 -8
rect 6 -20 10 -19
<< ntransistor >>
rect 7 -12 9 -8
<< ptransistor >>
rect -1 2 1 6
<< polycontact >>
rect -2 9 2 13
rect 6 -19 10 -15
<< ndcontact >>
rect 2 -12 6 -8
rect 10 -12 14 -8
<< pdcontact >>
rect -6 2 -2 6
rect 2 2 6 6
<< m2contact >>
rect -2 14 2 18
rect 6 -24 10 -20
<< end >>
