magic
tech scmos
timestamp 1385973147
<< metal1 >>
rect 94 62 135 66
rect -34 4 2 8
rect -34 -59 -30 4
rect 131 -1 135 62
rect 94 -5 135 -1
rect -34 -63 0 -59
rect -34 -127 -30 -63
rect 131 -69 135 -5
rect 93 -73 135 -69
rect -34 -131 1 -127
rect -34 -196 -30 -131
rect 131 -138 135 -73
rect 97 -142 135 -138
rect -34 -200 0 -196
rect -34 -265 -30 -200
rect 131 -207 135 -142
rect 95 -211 135 -207
rect -34 -269 0 -265
rect -34 -333 -30 -269
rect 131 -275 135 -211
rect 94 -279 135 -275
rect -34 -337 0 -333
rect -34 -400 -30 -337
rect 131 -342 135 -279
rect 96 -346 135 -342
rect -34 -404 0 -400
rect -34 -469 -30 -404
rect 131 -411 135 -346
rect 95 -415 135 -411
rect -34 -473 2 -469
rect -34 -538 -30 -473
rect 131 -480 135 -415
rect 97 -484 135 -480
rect -34 -542 2 -538
rect -34 -607 -30 -542
rect 131 -549 135 -484
rect 97 -553 135 -549
rect -34 -611 0 -607
rect -34 -676 -30 -611
rect 131 -618 135 -553
rect 92 -622 135 -618
rect -34 -680 4 -676
rect -34 -744 -30 -680
rect 131 -686 135 -622
rect 95 -690 135 -686
rect -34 -748 0 -744
rect -34 -813 -30 -748
rect 131 -755 135 -690
rect 93 -759 135 -755
rect -34 -817 0 -813
rect -34 -881 -30 -817
rect 131 -823 135 -759
rect 95 -827 135 -823
rect -34 -885 0 -881
rect -34 -950 -30 -885
rect 131 -892 135 -827
rect 94 -896 135 -892
rect -34 -954 0 -950
rect -34 -1019 -30 -954
rect 131 -961 135 -896
rect 96 -965 135 -961
rect -34 -1023 1 -1019
rect -34 -1087 -30 -1023
rect 131 -1029 135 -965
rect 95 -1033 135 -1029
rect -34 -1091 0 -1087
rect -34 -1154 -30 -1091
rect 131 -1096 135 -1033
rect 96 -1100 135 -1096
rect 131 -1101 135 -1100
rect -35 -1158 4 -1154
rect -34 -1159 -30 -1158
<< metal2 >>
rect 96 39 113 43
rect -17 31 0 35
rect -17 -32 -13 31
rect 109 -24 113 39
rect 94 -28 113 -24
rect -17 -36 2 -32
rect -17 -100 -13 -36
rect 109 -92 113 -28
rect 97 -96 113 -92
rect -17 -104 3 -100
rect -17 -169 -13 -104
rect 109 -161 113 -96
rect 94 -165 113 -161
rect -17 -173 0 -169
rect -17 -238 -13 -173
rect 109 -230 113 -165
rect 96 -234 113 -230
rect -17 -242 3 -238
rect -17 -306 -13 -242
rect 109 -298 113 -234
rect 97 -302 113 -298
rect -17 -310 2 -306
rect -17 -373 -13 -310
rect 109 -365 113 -302
rect 96 -369 113 -365
rect -17 -377 1 -373
rect -17 -442 -13 -377
rect 109 -434 113 -369
rect 95 -438 113 -434
rect -17 -446 4 -442
rect -17 -511 -13 -446
rect 109 -503 113 -438
rect 92 -507 113 -503
rect -17 -515 1 -511
rect -17 -580 -13 -515
rect 109 -572 113 -507
rect 96 -576 113 -572
rect -17 -584 0 -580
rect -17 -649 -13 -584
rect 109 -641 113 -576
rect 95 -645 114 -641
rect -17 -653 1 -649
rect -17 -717 -13 -653
rect 109 -709 113 -645
rect 95 -713 113 -709
rect -17 -721 1 -717
rect -17 -786 -13 -721
rect 109 -778 113 -713
rect 97 -782 113 -778
rect -17 -790 0 -786
rect -17 -854 -13 -790
rect 109 -846 113 -782
rect 97 -850 113 -846
rect -17 -858 0 -854
rect -17 -923 -13 -858
rect 109 -915 113 -850
rect 97 -919 113 -915
rect -17 -927 1 -923
rect -17 -992 -13 -927
rect 109 -984 113 -919
rect 96 -988 113 -984
rect -17 -996 0 -992
rect -17 -1060 -13 -996
rect 109 -1052 113 -988
rect 97 -1056 113 -1052
rect -17 -1064 3 -1060
rect -17 -1127 -13 -1064
rect 109 -1118 113 -1056
rect 105 -1119 113 -1118
rect 95 -1123 113 -1119
rect -17 -1131 2 -1127
use reg1  reg1_0
timestamp 1384799288
transform 1 0 20 0 1 62
box -20 -62 77 8
use reg1  reg1_1
timestamp 1384799288
transform 1 0 20 0 1 -5
box -20 -62 77 8
use reg1  reg1_2
timestamp 1384799288
transform 1 0 20 0 1 -73
box -20 -62 77 8
use reg1  reg1_3
timestamp 1384799288
transform 1 0 20 0 1 -142
box -20 -62 77 8
use reg1  reg1_4
timestamp 1384799288
transform 1 0 20 0 1 -211
box -20 -62 77 8
use reg1  reg1_5
timestamp 1384799288
transform 1 0 20 0 1 -279
box -20 -62 77 8
use reg1  reg1_6
timestamp 1384799288
transform 1 0 20 0 1 -346
box -20 -62 77 8
use reg1  reg1_7
timestamp 1384799288
transform 1 0 20 0 1 -415
box -20 -62 77 8
use reg1  reg1_8
timestamp 1384799288
transform 1 0 20 0 1 -484
box -20 -62 77 8
use reg1  reg1_9
timestamp 1384799288
transform 1 0 20 0 1 -553
box -20 -62 77 8
use reg1  reg1_10
timestamp 1384799288
transform 1 0 20 0 1 -622
box -20 -62 77 8
use reg1  reg1_11
timestamp 1384799288
transform 1 0 20 0 1 -690
box -20 -62 77 8
use reg1  reg1_12
timestamp 1384799288
transform 1 0 20 0 1 -759
box -20 -62 77 8
use reg1  reg1_13
timestamp 1384799288
transform 1 0 20 0 1 -827
box -20 -62 77 8
use reg1  reg1_14
timestamp 1384799288
transform 1 0 20 0 1 -896
box -20 -62 77 8
use reg1  reg1_15
timestamp 1384799288
transform 1 0 20 0 1 -965
box -20 -62 77 8
use reg1  reg1_16
timestamp 1384799288
transform 1 0 20 0 1 -1033
box -20 -62 77 8
use reg1  reg1_17
timestamp 1384799288
transform 1 0 20 0 1 -1100
box -20 -62 77 8
<< end >>
