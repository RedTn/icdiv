magic
tech scmos
timestamp 1384924723
<< pwell >>
rect -18 -31 13 -1
rect 201 -31 229 -12
rect 238 -31 472 2
<< nwell >>
rect -18 -1 13 31
rect 201 12 229 31
rect 238 2 472 31
<< polysilicon >>
rect 355 20 365 22
rect 392 22 416 25
rect -13 18 -11 20
rect 206 18 208 20
rect 222 18 224 20
rect 243 18 245 20
rect 250 18 252 20
rect 267 18 269 20
rect 283 18 285 20
rect 299 18 301 20
rect 307 18 309 20
rect 323 18 325 20
rect 331 18 333 20
rect 347 18 349 20
rect -13 3 -11 14
rect -14 -1 -11 3
rect -13 -14 -11 -1
rect 206 -14 208 14
rect 222 0 224 14
rect 243 11 245 14
rect 250 13 252 14
rect 250 11 253 13
rect 241 9 245 11
rect 241 5 243 9
rect 251 5 253 11
rect 239 1 243 5
rect 250 1 253 5
rect 267 4 269 14
rect 283 5 285 14
rect 299 5 301 14
rect 307 5 309 14
rect 323 12 325 14
rect 318 10 325 12
rect 318 5 320 10
rect 222 -2 226 0
rect 224 -10 226 -2
rect 222 -12 226 -10
rect 241 -10 243 1
rect 241 -12 245 -10
rect 222 -14 224 -12
rect 243 -14 245 -12
rect 251 -14 253 1
rect 266 0 269 4
rect 282 1 285 5
rect 298 1 301 5
rect 308 1 309 5
rect 316 1 320 5
rect 267 -14 269 0
rect 283 -6 285 1
rect 283 -12 285 -10
rect 299 -14 301 1
rect 307 -14 309 1
rect 318 -10 320 1
rect 318 -12 325 -10
rect 323 -14 325 -12
rect 331 -14 333 14
rect 347 -3 349 14
rect 355 5 357 20
rect 363 18 365 20
rect 371 18 373 20
rect 379 18 381 20
rect 395 18 397 20
rect 399 18 401 20
rect 407 18 409 20
rect 411 18 413 20
rect 428 18 430 20
rect 441 18 443 21
rect 457 18 459 20
rect 363 12 365 14
rect 371 5 373 14
rect 379 5 381 14
rect 395 13 397 14
rect 355 2 358 5
rect 370 2 373 5
rect 380 1 381 5
rect 346 -7 349 -3
rect 347 -14 349 -7
rect 359 -10 361 1
rect 367 -10 369 1
rect 359 -12 365 -10
rect 367 -12 373 -10
rect 363 -14 365 -12
rect 371 -14 373 -12
rect 379 -14 381 1
rect 388 11 397 13
rect 388 -5 390 11
rect 399 8 401 14
rect 407 13 409 14
rect 395 6 401 8
rect 404 11 409 13
rect 411 13 413 14
rect 411 11 416 13
rect 404 7 406 11
rect 414 10 416 11
rect 414 8 423 10
rect 420 7 423 8
rect 428 7 430 14
rect 441 11 443 14
rect 441 9 447 11
rect 444 7 447 9
rect 395 5 398 6
rect 395 0 398 1
rect 404 3 407 7
rect 428 3 431 7
rect 395 -2 402 0
rect 388 -9 391 -5
rect 388 -16 390 -9
rect 400 -15 402 -2
rect 404 -3 406 3
rect 420 -2 422 3
rect 404 -5 413 -3
rect 411 -11 413 -5
rect 419 -4 422 -2
rect 419 -11 421 -4
rect 428 -11 430 3
rect 444 0 447 3
rect 445 -9 447 0
rect 457 -6 459 14
rect 454 -8 459 -6
rect 427 -13 430 -11
rect 435 -11 447 -9
rect 388 -18 397 -16
rect 400 -17 405 -15
rect 411 -17 413 -15
rect 419 -17 421 -15
rect -13 -20 -11 -18
rect 206 -20 208 -18
rect 222 -20 224 -18
rect 243 -20 245 -18
rect 251 -20 253 -18
rect 267 -20 269 -18
rect 299 -20 301 -18
rect 307 -20 309 -18
rect 323 -20 325 -18
rect 331 -20 333 -18
rect 347 -20 349 -18
rect 363 -20 365 -18
rect 371 -20 373 -18
rect 379 -20 381 -18
rect 395 -19 397 -18
rect 403 -19 405 -17
rect 427 -19 429 -13
rect 435 -19 437 -11
rect 457 -14 459 -8
rect 457 -20 459 -18
rect 395 -25 397 -23
rect 403 -25 405 -23
rect 427 -25 429 -23
rect 435 -25 437 -23
<< ndiffusion >>
rect 282 -10 283 -6
rect 285 -10 286 -6
rect -14 -18 -13 -14
rect -11 -18 -10 -14
rect 205 -18 206 -14
rect 208 -18 209 -14
rect 221 -18 222 -14
rect 224 -18 225 -14
rect 242 -18 243 -14
rect 245 -18 246 -14
rect 250 -18 251 -14
rect 253 -18 254 -14
rect 266 -18 267 -14
rect 269 -18 270 -14
rect 298 -18 299 -14
rect 301 -18 302 -14
rect 306 -18 307 -14
rect 309 -18 310 -14
rect 322 -18 323 -14
rect 325 -18 331 -14
rect 333 -18 334 -14
rect 346 -18 347 -14
rect 349 -18 350 -14
rect 362 -18 363 -14
rect 365 -18 366 -14
rect 370 -18 371 -14
rect 373 -18 374 -14
rect 378 -18 379 -14
rect 381 -18 382 -14
rect 410 -15 411 -11
rect 413 -15 414 -11
rect 418 -15 419 -11
rect 421 -15 422 -11
rect 456 -18 457 -14
rect 459 -18 460 -14
rect 394 -23 395 -19
rect 397 -23 398 -19
rect 402 -23 403 -19
rect 405 -23 406 -19
rect 426 -23 427 -19
rect 429 -23 430 -19
rect 434 -23 435 -19
rect 437 -23 438 -19
<< pdiffusion >>
rect -14 14 -13 18
rect -11 14 -10 18
rect 205 14 206 18
rect 208 14 209 18
rect 221 14 222 18
rect 224 14 225 18
rect 242 14 243 18
rect 245 14 250 18
rect 252 14 254 18
rect 266 14 267 18
rect 269 14 270 18
rect 282 14 283 18
rect 285 14 286 18
rect 290 14 299 18
rect 301 14 307 18
rect 309 14 310 18
rect 322 14 323 18
rect 325 14 326 18
rect 330 14 331 18
rect 333 14 334 18
rect 346 14 347 18
rect 349 14 350 18
rect 362 14 363 18
rect 365 14 371 18
rect 373 14 379 18
rect 381 14 382 18
rect 394 14 395 18
rect 397 14 399 18
rect 401 14 402 18
rect 406 14 407 18
rect 409 14 411 18
rect 413 14 414 18
rect 426 14 428 18
rect 430 14 441 18
rect 443 14 444 18
rect 456 14 457 18
rect 459 14 460 18
<< metal1 >>
rect 178 128 209 132
rect 155 109 197 113
rect 225 109 422 113
rect -19 102 174 106
rect -101 83 54 87
rect 58 83 166 87
rect 191 83 383 87
rect -60 73 151 77
rect 290 75 449 79
rect 378 67 391 71
rect 395 67 415 71
rect 419 67 439 71
rect 193 59 235 63
rect 239 59 358 63
rect 193 39 197 59
rect 207 51 243 55
rect 247 51 278 55
rect 282 51 324 55
rect 328 51 431 55
rect 215 43 294 47
rect 298 43 310 47
rect 314 43 407 47
rect 144 35 193 39
rect 231 35 302 39
rect 306 35 342 39
rect 346 35 366 39
rect -18 27 -10 31
rect 0 27 8 31
rect 199 27 217 31
rect 221 27 238 31
rect -84 15 -27 19
rect -18 18 -14 27
rect -10 8 -6 14
rect -73 -27 -69 0
rect -32 -27 -28 0
rect -19 -1 -18 3
rect -10 -14 -6 4
rect 1 0 5 14
rect 98 -17 102 15
rect 194 4 198 16
rect 201 18 205 27
rect 217 18 221 27
rect 242 27 262 31
rect 238 18 242 24
rect 266 27 278 31
rect 262 18 266 24
rect 282 27 318 31
rect 278 18 282 24
rect 310 18 314 27
rect 322 27 342 31
rect 318 18 322 24
rect 334 18 338 27
rect 346 27 358 31
rect 342 18 346 24
rect 362 28 431 31
rect 362 27 385 28
rect 395 27 413 28
rect 423 27 431 28
rect 448 27 460 31
rect 464 27 468 31
rect 358 18 362 24
rect 392 21 393 24
rect 390 18 394 21
rect 402 18 406 27
rect 416 18 420 21
rect 423 18 426 19
rect 418 14 422 18
rect 444 18 448 27
rect 452 18 456 27
rect 209 4 213 14
rect 225 4 229 14
rect 235 5 239 6
rect 194 0 202 4
rect 209 0 211 4
rect 209 -14 213 0
rect 218 -4 222 0
rect 225 0 227 4
rect 246 5 250 6
rect 254 4 258 14
rect 270 5 274 14
rect 270 4 278 5
rect 258 0 262 4
rect 274 1 278 4
rect 286 2 290 14
rect 225 -14 229 0
rect 254 -2 258 0
rect 246 -6 258 -2
rect 246 -14 250 -6
rect 270 -14 274 0
rect 294 5 298 6
rect 306 6 307 8
rect 302 5 307 6
rect 312 5 316 6
rect 286 -6 290 -2
rect 326 -3 330 14
rect 334 5 338 6
rect 350 -3 354 14
rect 382 12 386 14
rect 382 10 387 12
rect 358 5 362 6
rect 366 5 370 6
rect 382 8 383 10
rect 374 5 378 6
rect 431 7 435 8
rect 374 1 376 5
rect -18 -27 -14 -18
rect 201 -27 205 -18
rect 217 -27 221 -18
rect 238 -24 242 -18
rect -73 -31 -10 -27
rect 0 -31 6 -27
rect 199 -31 217 -27
rect 221 -31 238 -27
rect 254 -27 258 -18
rect 294 -10 314 -6
rect 330 -7 342 -3
rect 383 -6 387 6
rect 398 1 399 5
rect 419 3 420 7
rect 443 3 444 7
rect 407 2 411 3
rect 460 0 464 14
rect 414 -3 442 0
rect 278 -14 282 -10
rect 294 -14 298 -10
rect 310 -14 314 -10
rect 334 -14 338 -7
rect 350 -14 354 -7
rect 366 -10 387 -6
rect 391 -10 395 -9
rect 366 -14 370 -10
rect 382 -14 386 -10
rect 406 -11 410 -10
rect 278 -18 294 -14
rect 398 -15 406 -11
rect 414 -11 418 -3
rect 422 -11 426 -10
rect 262 -24 266 -18
rect 242 -31 262 -27
rect 302 -24 306 -18
rect 266 -31 302 -27
rect 318 -24 322 -18
rect 306 -31 318 -27
rect 342 -24 346 -18
rect 322 -31 342 -27
rect 358 -27 362 -18
rect 374 -24 378 -18
rect 398 -19 402 -15
rect 414 -19 418 -15
rect 430 -19 434 -18
rect 346 -31 374 -27
rect 414 -23 422 -19
rect 438 -19 442 -3
rect 449 -5 453 -4
rect 460 -14 464 -4
rect 390 -27 394 -23
rect 406 -27 410 -23
rect 452 -27 456 -18
rect 378 -31 397 -27
rect 435 -31 452 -27
rect 456 -31 460 -27
rect 464 -31 472 -27
rect 282 -39 294 -35
<< metal2 >>
rect -23 106 -19 122
rect -105 0 -101 83
rect -64 0 -60 73
rect -23 3 -19 102
rect 1 18 5 110
rect 54 35 58 83
rect 151 77 155 109
rect 174 106 178 128
rect 98 35 140 39
rect 151 35 155 73
rect 213 68 217 93
rect 182 64 217 68
rect 98 19 102 35
rect 182 8 186 64
rect 193 25 197 35
rect 193 21 198 25
rect 194 20 198 21
rect -6 4 6 8
rect -10 -19 -6 4
rect -91 -23 -6 -19
rect 98 -31 102 -21
rect 203 -31 207 51
rect 211 4 215 43
rect 227 4 231 35
rect 235 10 239 59
rect 243 10 247 51
rect 243 6 246 10
rect 218 -31 222 -8
rect 58 -35 102 -31
rect 155 -35 222 -31
rect 254 -34 258 0
rect 270 -34 274 0
rect 246 -38 258 -34
rect 246 -42 250 -38
rect 254 -42 258 -38
rect 262 -38 274 -34
rect 262 -42 266 -38
rect 270 -42 274 -38
rect 278 -35 282 51
rect 278 -42 282 -39
rect 286 2 290 75
rect 294 10 298 43
rect 302 10 306 35
rect 310 10 314 43
rect 324 24 328 51
rect 324 20 338 24
rect 334 10 338 20
rect 310 6 312 10
rect 286 -42 290 -2
rect 294 -42 298 -39
rect 326 -42 330 -7
rect 342 -42 346 35
rect 358 10 362 59
rect 366 10 370 35
rect 374 10 378 67
rect 383 10 387 83
rect 422 77 426 109
rect 350 -42 354 -7
rect 391 -10 395 67
rect 407 2 411 43
rect 415 7 418 67
rect 423 63 426 77
rect 422 23 426 63
rect 422 12 426 19
rect 423 11 426 12
rect 431 12 435 51
rect 399 -31 402 1
rect 423 2 427 11
rect 439 7 443 67
rect 423 -2 434 2
rect 410 -10 422 -6
rect 430 -14 434 -2
rect 449 0 453 75
rect 399 -42 403 -31
rect 452 -42 456 -31
rect 460 -42 464 -4
rect 468 -42 472 27
<< ntransistor >>
rect 283 -10 285 -6
rect -13 -18 -11 -14
rect 206 -18 208 -14
rect 222 -18 224 -14
rect 243 -18 245 -14
rect 251 -18 253 -14
rect 267 -18 269 -14
rect 299 -18 301 -14
rect 307 -18 309 -14
rect 323 -18 325 -14
rect 331 -18 333 -14
rect 347 -18 349 -14
rect 363 -18 365 -14
rect 371 -18 373 -14
rect 379 -18 381 -14
rect 411 -15 413 -11
rect 419 -15 421 -11
rect 457 -18 459 -14
rect 395 -23 397 -19
rect 403 -23 405 -19
rect 427 -23 429 -19
rect 435 -23 437 -19
<< ptransistor >>
rect -13 14 -11 18
rect 206 14 208 18
rect 222 14 224 18
rect 243 14 245 18
rect 250 14 252 18
rect 267 14 269 18
rect 283 14 285 18
rect 299 14 301 18
rect 307 14 309 18
rect 323 14 325 18
rect 331 14 333 18
rect 347 14 349 18
rect 363 14 365 18
rect 371 14 373 18
rect 379 14 381 18
rect 395 14 397 18
rect 399 14 401 18
rect 407 14 409 18
rect 411 14 413 18
rect 428 14 430 18
rect 441 14 443 18
rect 457 14 459 18
<< polycontact >>
rect 388 21 392 25
rect 416 21 420 25
rect -18 -1 -14 3
rect 202 0 206 4
rect 218 0 222 4
rect 235 1 239 5
rect 246 1 250 5
rect 262 0 266 4
rect 278 1 282 5
rect 294 1 298 5
rect 304 1 308 5
rect 312 1 316 5
rect 333 1 337 5
rect 358 1 362 5
rect 366 1 370 5
rect 376 1 380 5
rect 342 -7 346 -3
rect 394 1 398 5
rect 407 3 411 7
rect 420 3 424 7
rect 431 3 435 7
rect 444 3 448 7
rect 391 -9 395 -5
rect 450 -9 454 -5
<< ndcontact >>
rect 278 -10 282 -6
rect 286 -10 290 -6
rect -18 -18 -14 -14
rect -10 -18 -6 -14
rect 201 -18 205 -14
rect 209 -18 213 -14
rect 217 -18 221 -14
rect 225 -18 229 -14
rect 238 -18 242 -14
rect 246 -18 250 -14
rect 254 -18 258 -14
rect 262 -18 266 -14
rect 270 -18 274 -14
rect 294 -18 298 -14
rect 302 -18 306 -14
rect 310 -18 314 -14
rect 318 -18 322 -14
rect 334 -18 338 -14
rect 342 -18 346 -14
rect 350 -18 354 -14
rect 358 -18 362 -14
rect 366 -18 370 -14
rect 374 -18 378 -14
rect 382 -18 386 -14
rect 406 -15 410 -11
rect 414 -15 418 -11
rect 422 -15 426 -11
rect 452 -18 456 -14
rect 460 -18 464 -14
rect 390 -23 394 -19
rect 398 -23 402 -19
rect 406 -23 410 -19
rect 422 -23 426 -19
rect 430 -23 434 -19
rect 438 -23 442 -19
<< pdcontact >>
rect -18 14 -14 18
rect -10 14 -6 18
rect 201 14 205 18
rect 209 14 213 18
rect 217 14 221 18
rect 225 14 229 18
rect 238 14 242 18
rect 254 14 258 18
rect 262 14 266 18
rect 270 14 274 18
rect 278 14 282 18
rect 286 14 290 18
rect 310 14 314 18
rect 318 14 322 18
rect 326 14 330 18
rect 334 14 338 18
rect 342 14 346 18
rect 350 14 354 18
rect 358 14 362 18
rect 382 14 386 18
rect 390 14 394 18
rect 402 14 406 18
rect 414 14 418 18
rect 422 14 426 18
rect 444 14 448 18
rect 452 14 456 18
rect 460 14 464 18
<< m2contact >>
rect 174 128 178 132
rect 1 110 5 114
rect 151 109 155 113
rect 422 109 426 113
rect -23 102 -19 106
rect -105 83 -101 87
rect 54 83 58 87
rect 383 83 387 87
rect -64 73 -60 77
rect 151 73 155 77
rect 286 75 290 79
rect 449 75 453 79
rect 374 67 378 71
rect 391 67 395 71
rect 415 67 419 71
rect 439 67 443 71
rect 235 59 239 63
rect 358 59 362 63
rect 203 51 207 55
rect 243 51 247 55
rect 278 51 282 55
rect 324 51 328 55
rect 431 51 435 55
rect 211 43 215 47
rect 294 43 298 47
rect 310 43 314 47
rect 407 43 411 47
rect 140 35 144 39
rect 193 35 197 39
rect 227 35 231 39
rect 302 35 306 39
rect 342 35 346 39
rect 366 35 370 39
rect -27 15 -23 19
rect -10 4 -6 8
rect -105 -4 -101 0
rect -64 -4 -60 0
rect -23 -1 -19 3
rect 1 14 5 18
rect 1 -4 5 0
rect 98 15 102 19
rect 194 16 198 20
rect 468 27 472 31
rect 423 19 427 23
rect 235 6 239 10
rect 211 0 215 4
rect 218 -8 222 -4
rect 227 0 231 4
rect 246 6 250 10
rect 254 0 258 4
rect 270 0 274 4
rect 286 -2 290 2
rect 294 6 298 10
rect 302 6 306 10
rect 312 6 316 10
rect 334 6 338 10
rect 358 6 362 10
rect 366 6 370 10
rect 374 6 378 10
rect 383 6 387 10
rect 431 8 435 12
rect 98 -21 102 -17
rect 326 -7 330 -3
rect 350 -7 354 -3
rect 399 1 403 5
rect 415 3 419 7
rect 439 3 443 7
rect 407 -2 411 2
rect 391 -14 395 -10
rect 406 -10 410 -6
rect 422 -10 426 -6
rect 430 -18 434 -14
rect 449 -4 453 0
rect 460 -4 464 0
rect 452 -31 456 -27
rect 278 -39 282 -35
rect 294 -39 298 -35
<< psubstratepcontact >>
rect -10 -31 0 -27
rect 217 -31 221 -27
rect 238 -31 242 -24
rect 262 -31 266 -24
rect 302 -31 306 -24
rect 318 -31 322 -24
rect 342 -31 346 -24
rect 374 -31 378 -24
rect 397 -31 435 -27
rect 460 -31 464 -27
<< nsubstratencontact >>
rect -10 27 0 31
rect 217 27 221 31
rect 238 24 242 31
rect 262 24 266 31
rect 278 24 282 31
rect 318 24 322 31
rect 342 24 346 31
rect 358 24 362 31
rect 431 27 448 31
rect 460 27 464 31
use transgate  transgate_0
timestamp 1384720590
transform 1 0 176 0 1 88
box -10 -24 18 18
use transgate  transgate_1
timestamp 1384720590
transform 1 0 207 0 1 114
box -10 -24 18 18
use transgate  transgate_3
timestamp 1384720590
transform 1 0 -91 0 -1 -5
box -10 -24 18 18
use transgate  transgate_2
timestamp 1384720590
transform 1 0 -50 0 -1 -5
box -10 -24 18 18
use dflipflop  dflipflop_0
timestamp 1384718467
transform 1 0 25 0 1 27
box -20 -62 77 8
use dflipflop  dflipflop_1
timestamp 1384718467
transform 1 0 122 0 1 27
box -20 -62 77 8
<< labels >>
rlabel metal2 270 -42 274 0 5 loadb
rlabel metal2 254 -42 258 0 5 load
rlabel metal2 286 -42 290 -38 5 sel1
rlabel metal2 326 -42 330 -7 5 shift
rlabel metal2 350 -42 354 -7 5 shiftb
rlabel m2contact 374 67 378 71 1 start
rlabel m2contact 383 83 387 87 1 xout
rlabel metal1 197 59 235 63 1 x
rlabel metal1 207 51 243 55 1 y
rlabel m2contact 422 109 426 113 1 yout
rlabel metal2 182 8 186 68 7 resetb
rlabel metal2 54 35 58 83 7 xin
rlabel metal2 151 35 155 73 7 yin
rlabel metal2 262 -42 266 -34 5 sel0
rlabel metal2 278 -42 282 51 5 inbit
rlabel metal2 342 -42 346 35 5 add
rlabel m2contact 1 110 5 114 7 Clk
rlabel metal2 -23 106 -19 122 1 reset
rlabel metal2 399 -42 403 -31 5 sign
rlabel metal2 460 -42 464 -4 5 sel1b
rlabel metal2 468 -42 472 27 5 Vdd
rlabel metal2 452 -42 456 -31 5 Gnd
rlabel metal2 246 -42 250 -34 5 sel0b
rlabel metal2 294 -42 298 -39 5 addb
<< end >>
