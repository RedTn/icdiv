magic
tech scmos
timestamp 1385529037
<< metal1 >>
rect -29 220 108 224
rect 117 220 341 224
rect -29 206 119 210
rect 128 206 341 210
rect -29 188 255 192
rect 263 188 341 192
rect -29 173 266 177
rect 273 173 341 177
rect 62 158 211 164
rect 216 157 281 164
rect 216 156 289 157
rect -29 135 55 139
rect 237 137 341 141
rect 182 -28 201 -24
rect 182 -29 207 -28
rect 182 -31 185 -29
rect -29 -37 162 -33
rect 235 -37 341 -33
rect -29 -49 155 -45
rect 240 -49 341 -45
rect -29 -57 155 -53
rect 240 -57 341 -53
rect -29 -86 155 -82
rect 240 -86 341 -82
rect -11 -91 155 -90
rect -29 -94 155 -91
rect 240 -94 341 -90
rect -29 -95 79 -94
rect 182 -130 186 -103
rect 3 -143 145 -139
rect -29 -166 143 -162
rect 240 -166 341 -162
rect -29 -174 143 -170
rect 240 -174 341 -170
rect -29 -200 14 -196
rect 25 -197 79 -196
rect 25 -201 147 -197
rect 236 -201 341 -197
rect 191 -214 192 -210
rect 196 -214 280 -210
rect 290 -214 292 -210
<< metal2 >>
rect 58 146 62 158
rect 66 150 71 319
rect 109 148 115 219
rect 119 147 125 205
rect 254 185 255 192
rect 254 174 261 185
rect 211 146 216 155
rect 255 143 260 174
rect 266 143 271 173
rect -4 -137 3 73
rect 17 -195 24 11
rect 201 -24 207 -4
rect 201 -29 207 -28
rect 181 -135 182 -131
rect 187 -135 196 -131
rect 192 -136 196 -135
rect 192 -210 196 -200
rect 281 -209 289 157
<< m2contact >>
rect 108 219 117 228
rect 119 205 128 211
rect 255 185 263 194
rect 266 173 273 178
rect 58 158 62 165
rect 211 155 216 164
rect 281 157 289 164
rect 16 11 24 15
rect 201 -28 208 -24
rect 155 -49 159 -45
rect 236 -49 240 -45
rect 155 -57 159 -53
rect 236 -57 240 -53
rect 155 -86 159 -82
rect 236 -86 240 -82
rect 155 -94 159 -90
rect 236 -94 240 -90
rect 182 -136 187 -130
rect -5 -145 3 -137
rect 143 -166 147 -162
rect 236 -166 240 -162
rect 143 -174 147 -170
rect 236 -174 240 -170
rect 14 -203 25 -195
rect 192 -214 196 -210
rect 280 -216 290 -209
use real31mux  real31mux_0
timestamp 1385529037
transform 1 0 -9 0 1 7
box 6 -14 280 146
use shiftv2  shiftv2_0
timestamp 1385333955
transform 1 0 190 0 1 -102
box -35 -8 50 73
use dflipfloplabels  dflipfloplabels_0
timestamp 1384799288
transform 1 0 163 0 1 -143
box -20 -62 77 8
<< end >>
