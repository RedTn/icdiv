magic
tech scmos
timestamp 1385343589
<< pwell >>
rect -50 -34 36 -8
rect -51 -109 35 -68
rect -62 -172 37 -145
rect -67 -223 37 -197
<< nwell >>
rect -42 -5 32 25
rect -47 -67 32 -37
rect -47 -140 36 -110
rect -74 -193 36 -175
<< polysilicon >>
rect -14 19 -11 22
rect -27 -56 -24 -17
rect -14 -18 -11 16
rect -3 12 0 22
rect 7 19 10 21
rect -3 4 0 9
rect 7 4 10 16
rect -3 -10 0 1
rect 7 -10 10 1
rect -14 -41 -11 -21
rect -3 -27 0 -13
rect 7 -18 10 -13
rect 7 -22 10 -21
rect 7 -26 8 -22
rect -3 -41 0 -30
rect 9 -41 12 -36
rect -14 -56 -11 -44
rect -3 -48 0 -44
rect -27 -83 -24 -59
rect -14 -75 -11 -59
rect -3 -75 0 -51
rect 9 -60 12 -44
rect 9 -75 12 -63
rect -14 -83 -11 -78
rect -27 -91 -24 -86
rect -27 -127 -24 -108
rect -14 -127 -11 -86
rect -3 -91 0 -78
rect -3 -117 0 -94
rect 9 -99 12 -78
rect 9 -104 12 -102
rect -53 -161 -47 -158
rect -53 -177 -50 -161
rect -27 -157 -24 -130
rect -14 -136 -11 -130
rect -3 -136 0 -120
rect -14 -150 -11 -139
rect -3 -150 0 -139
rect -14 -157 -11 -153
rect -53 -218 -50 -180
rect -40 -178 -37 -160
rect -27 -162 -24 -160
rect -14 -162 -11 -160
rect -3 -166 0 -153
rect -3 -171 0 -169
rect -33 -173 -29 -172
rect -33 -176 3 -173
rect -40 -181 -26 -178
rect 0 -179 3 -176
rect -29 -186 -26 -181
rect -29 -210 -26 -189
rect 0 -199 3 -182
rect 0 -204 3 -202
rect -29 -215 -26 -213
rect -53 -223 -50 -221
<< ndiffusion >>
rect -5 -13 -3 -10
rect 0 -13 7 -10
rect 10 -13 24 -10
rect -15 -21 -14 -18
rect -11 -21 -9 -18
rect 5 -21 7 -18
rect 10 -21 24 -18
rect -5 -30 -3 -27
rect 0 -30 24 -27
rect -17 -78 -14 -75
rect -11 -78 -3 -75
rect 0 -78 9 -75
rect 12 -78 13 -75
rect -29 -86 -27 -83
rect -24 -86 -22 -83
rect -18 -86 -14 -83
rect -11 -86 -10 -83
rect -6 -94 -3 -91
rect 0 -94 1 -91
rect 5 -102 9 -99
rect 12 -102 13 -99
rect -15 -153 -14 -150
rect -11 -153 -3 -150
rect 0 -153 2 -150
rect -29 -160 -27 -157
rect -24 -160 -23 -157
rect -19 -160 -14 -157
rect -11 -160 -10 -157
rect -19 -169 -3 -166
rect 0 -169 2 -166
rect -5 -202 0 -199
rect 3 -202 10 -199
rect -31 -213 -29 -210
rect -26 -213 10 -210
rect -56 -221 -53 -218
rect -50 -221 10 -218
<< pdiffusion >>
rect -16 16 -14 19
rect -11 16 -9 19
rect 5 16 7 19
rect 10 16 11 19
rect -5 9 -3 12
rect 0 9 2 12
rect -5 1 -3 4
rect 0 1 7 4
rect 10 1 11 4
rect -16 -44 -14 -41
rect -11 -44 -3 -41
rect 0 -44 9 -41
rect 12 -44 13 -41
rect -28 -59 -27 -56
rect -24 -59 -21 -56
rect -5 -51 -3 -48
rect 0 -51 1 -48
rect -17 -59 -14 -56
rect -11 -59 -9 -56
rect 8 -63 9 -60
rect 12 -63 13 -60
rect -4 -120 -3 -117
rect 0 -120 17 -117
rect -28 -130 -27 -127
rect -24 -130 -19 -127
rect -15 -130 -14 -127
rect -11 -130 -9 -127
rect -15 -139 -14 -136
rect -11 -139 -3 -136
rect 0 -139 1 -136
rect -56 -180 -53 -177
rect -50 -180 -46 -177
rect -5 -182 0 -179
rect 3 -182 5 -179
rect -31 -189 -29 -186
rect -26 -189 -20 -186
<< metal1 >>
rect -5 16 1 19
rect -20 11 -16 16
rect -8 12 -5 16
rect 12 12 15 16
rect 18 17 19 20
rect 18 12 21 17
rect -46 7 -16 11
rect 6 9 21 12
rect -46 -158 -43 7
rect -20 4 -16 7
rect 12 5 15 9
rect -20 1 -9 4
rect -20 -3 -16 1
rect -19 -10 -16 -3
rect -19 -13 -9 -10
rect -23 -16 -16 -13
rect -19 -17 -16 -16
rect -5 -21 1 -18
rect -8 -26 -5 -22
rect 9 -32 12 -26
rect -33 -44 -20 -41
rect 18 -41 21 9
rect -32 -56 -28 -44
rect 24 1 27 12
rect 24 -8 32 1
rect 24 -9 36 -8
rect 24 -10 32 -9
rect 28 -12 32 -10
rect 24 -18 27 -14
rect 24 -27 27 -22
rect -20 -51 -9 -48
rect -20 -55 -17 -51
rect 1 -53 5 -52
rect 13 -49 17 -45
rect 13 -53 14 -49
rect -2 -55 17 -53
rect -32 -63 -28 -60
rect -40 -67 -28 -63
rect -8 -56 17 -55
rect -21 -64 -17 -59
rect -5 -58 1 -56
rect 14 -59 17 -56
rect 4 -64 8 -63
rect 13 -64 17 -63
rect -21 -67 8 -64
rect 14 -65 17 -64
rect -40 -156 -37 -67
rect -32 -75 -28 -67
rect 24 -75 27 -31
rect -32 -78 -21 -75
rect -32 -83 -29 -78
rect 17 -79 27 -75
rect 13 -83 17 -79
rect -6 -86 17 -83
rect -21 -91 -18 -87
rect 13 -91 17 -86
rect -21 -95 -10 -91
rect 5 -94 17 -91
rect -21 -99 -18 -95
rect 13 -99 17 -94
rect -21 -102 1 -99
rect 24 -87 27 -79
rect -34 -108 -29 -104
rect -34 -113 -30 -108
rect 4 -113 17 -110
rect 17 -117 21 -113
rect -19 -120 -8 -117
rect -19 -127 -15 -120
rect 17 -127 20 -121
rect -5 -130 9 -127
rect -32 -142 -29 -131
rect -19 -135 -16 -131
rect 13 -130 16 -127
rect 1 -142 5 -140
rect -32 -145 5 -142
rect -32 -150 -29 -145
rect -32 -153 -19 -150
rect -32 -156 -29 -153
rect 3 -155 6 -154
rect 24 -155 27 -94
rect 3 -156 27 -155
rect 3 -157 23 -156
rect -33 -168 -29 -160
rect -6 -158 23 -157
rect -6 -161 6 -158
rect -22 -165 -19 -161
rect 3 -165 6 -161
rect 16 -172 19 -165
rect -26 -175 19 -172
rect -19 -178 -16 -175
rect -42 -181 -16 -178
rect 16 -179 19 -175
rect -59 -218 -56 -181
rect -19 -185 -16 -181
rect 9 -182 19 -179
rect -35 -196 -32 -190
rect -8 -199 -5 -183
rect 16 -186 19 -182
rect 23 -199 27 -169
rect -35 -209 -32 -200
rect 14 -203 20 -199
rect 11 -204 20 -203
rect 11 -205 27 -204
rect 11 -209 14 -205
rect 11 -217 14 -213
<< metal2 >>
rect 18 -109 21 -65
rect -36 -117 -34 -113
rect -36 -196 -32 -117
rect 16 -161 19 -131
<< ntransistor >>
rect -3 -13 0 -10
rect 7 -13 10 -10
rect -14 -21 -11 -18
rect 7 -21 10 -18
rect -3 -30 0 -27
rect -14 -78 -11 -75
rect -3 -78 0 -75
rect 9 -78 12 -75
rect -27 -86 -24 -83
rect -14 -86 -11 -83
rect -3 -94 0 -91
rect 9 -102 12 -99
rect -14 -153 -11 -150
rect -3 -153 0 -150
rect -27 -160 -24 -157
rect -14 -160 -11 -157
rect -3 -169 0 -166
rect 0 -202 3 -199
rect -29 -213 -26 -210
rect -53 -221 -50 -218
<< ptransistor >>
rect -14 16 -11 19
rect 7 16 10 19
rect -3 9 0 12
rect -3 1 0 4
rect 7 1 10 4
rect -14 -44 -11 -41
rect -3 -44 0 -41
rect 9 -44 12 -41
rect -27 -59 -24 -56
rect -3 -51 0 -48
rect -14 -59 -11 -56
rect 9 -63 12 -60
rect -3 -120 0 -117
rect -27 -130 -24 -127
rect -14 -130 -11 -127
rect -14 -139 -11 -136
rect -3 -139 0 -136
rect -53 -180 -50 -177
rect 0 -182 3 -179
rect -29 -189 -26 -186
<< polycontact >>
rect -27 -17 -23 -13
rect 8 -26 12 -22
rect 8 -36 12 -32
rect -29 -108 -24 -104
rect -47 -162 -43 -158
rect -40 -160 -36 -156
rect -33 -172 -29 -168
<< ndcontact >>
rect -19 -21 -15 -17
rect -9 -14 -5 -10
rect -9 -22 -5 -18
rect -9 -30 -5 -26
rect 24 -14 28 -10
rect 1 -22 5 -18
rect 24 -22 28 -18
rect 24 -31 28 -27
rect -21 -79 -17 -75
rect -33 -87 -29 -83
rect -22 -87 -18 -83
rect -10 -87 -6 -83
rect -10 -95 -6 -91
rect 1 -95 5 -91
rect 13 -79 17 -75
rect 1 -103 5 -99
rect 13 -103 17 -99
rect -33 -160 -29 -156
rect -19 -153 -15 -149
rect -23 -161 -19 -157
rect -10 -161 -6 -157
rect -23 -169 -19 -165
rect 2 -154 6 -150
rect 2 -169 6 -165
rect -35 -213 -31 -209
rect -9 -203 -5 -199
rect 10 -203 14 -199
rect 10 -213 14 -209
rect -60 -222 -56 -218
rect 10 -221 14 -217
<< pdcontact >>
rect -20 16 -16 20
rect -9 16 -5 20
rect 1 16 5 20
rect 11 16 15 20
rect -9 8 -5 12
rect 2 8 6 12
rect -9 0 -5 4
rect 11 1 15 5
rect -20 -44 -16 -40
rect -32 -60 -28 -56
rect -21 -59 -17 -55
rect -9 -52 -5 -48
rect -9 -60 -5 -56
rect 1 -52 5 -48
rect 4 -63 8 -59
rect 13 -45 21 -41
rect 13 -63 17 -59
rect -8 -121 -4 -117
rect -32 -131 -28 -127
rect -19 -131 -15 -127
rect -19 -139 -15 -135
rect -9 -131 -5 -127
rect 17 -121 21 -117
rect 1 -140 5 -136
rect -60 -181 -56 -177
rect -46 -181 -42 -177
rect -9 -183 -5 -179
rect -35 -190 -31 -186
rect -20 -189 -16 -185
rect 5 -183 9 -179
<< m2contact >>
rect 14 -69 18 -65
rect 17 -113 21 -109
rect -34 -117 -30 -113
rect 16 -131 20 -127
rect 16 -165 20 -161
rect -36 -200 -32 -196
<< psubstratepcontact >>
rect 32 -14 36 -9
rect 24 -94 28 -87
rect 23 -169 31 -156
rect 20 -204 30 -199
<< nsubstratencontact >>
rect 19 17 23 21
rect 14 -53 20 -49
rect 9 -132 13 -127
rect 15 -191 19 -186
<< labels >>
rlabel metal1 -59 -200 -56 -197 1 a
rlabel metal1 -35 -200 -32 -192 1 b
rlabel metal1 -8 -194 -5 -190 1 c
rlabel polysilicon 7 13 10 16 1 ain
rlabel polysilicon -3 12 0 15 1 bin
rlabel polysilicon -14 12 -11 15 1 cin
rlabel metal1 -45 -33 -43 -30 1 aa
rlabel metal1 24 5 27 11 1 GND
rlabel metal1 18 5 21 10 1 Vdd
rlabel metal1 -40 -150 -37 -145 1 bb
rlabel metal1 -31 -149 -30 -145 1 cc
<< end >>
